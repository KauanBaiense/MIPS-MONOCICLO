memoriaMIPS_inst : memoriaMIPS PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
