package memReg is
    type Lista_registradores is array (31 downto 0) of STD_LOGIC_VECTOR(4 downto 0);
  end package memReg;
  
  package body memReg is
  end package body memReg;